magic
tech sky130A
magscale 1 2
timestamp 1742825900
<< locali >>
rect -1080 796 -888 1084
rect 72 796 264 1084
rect -1196 790 396 796
rect -1196 610 -690 790
rect -510 610 396 790
rect -1196 604 396 610
<< viali >>
rect -690 610 -510 790
<< metal1 >>
rect -312 4604 196 4796
rect -824 3894 -760 4250
rect -824 3171 -760 3459
rect -830 3107 -824 3171
rect -760 3107 -754 3171
rect -824 3022 -760 3107
rect -824 2311 -760 2650
rect -824 1520 -760 1836
rect -696 796 -504 4496
rect 4 3996 196 4604
rect -296 3804 196 3996
rect -212 3171 -148 3177
rect -212 3101 -148 3107
rect 4 2396 196 3804
rect -296 2204 196 2396
rect 4 1396 196 2204
rect -296 1204 196 1396
rect -702 790 -498 796
rect -702 610 -690 790
rect -510 610 -498 790
rect -702 604 -498 610
<< via1 >>
rect -824 3107 -760 3171
rect -212 3107 -148 3171
<< metal2 >>
rect -824 3171 -760 3177
rect -1100 3107 -824 3171
rect -760 3107 -212 3171
rect -148 3107 -142 3171
rect -824 3101 -760 3107
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ~/pro/aicex/ip/jnw_ex_sky130a/design/JNW_ATR_SKY130A
timestamp 1737385461
transform 1 0 -984 0 1 4076
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1737385461
transform 1 0 -984 0 1 884
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1737385461
transform 1 0 -984 0 1 1682
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1737385461
transform 1 0 -984 0 1 2480
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1737385461
transform 1 0 -984 0 1 3278
box -184 -128 1336 928
<< labels >>
flabel metal2 -1100 3107 -1036 3171 0 FreeSans 1600 0 0 0 IBPS_5U
port 1 nsew
flabel metal1 4 2838 196 3030 0 FreeSans 1600 0 0 0 IBNS_20U
port 3 nsew
flabel locali -1196 604 -1004 796 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
<< end >>
